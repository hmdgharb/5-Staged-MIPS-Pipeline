library verilog;
use verilog.vl_types.all;
entity bench is
end bench;
